module neon

pub enum KeyCode {
	unknown
	@return // 'return' is a reserved keyword
	escape
	backspace
	tab
	space
	exclaim
	dbl_apostrophe
	hash
	dollar
	percent
	ampersand
	apostrophe
	left_paren
	right_paren
	asterisk
	plus
	comma
	minus
	period
	slash
	num0
	num1
	num2
	num3
	num4
	num5
	num6
	num7
	num8
	num9
	colon
	semicolon
	less
	equals
	greater
	question
	at
	left_bracket
	backslash
	right_bracket
	caret
	underscore
	grave
	a
	b
	c
	d
	e
	f
	g
	h
	i
	j
	k
	l
	m
	n
	o
	p
	q
	r
	s
	t
	u
	v
	w
	x
	y
	z
	left_brace
	pipe
	right_brace
	tilde
	delete
	plus_minus
	caps_lock
	f1
	f2
	f3
	f4
	f5
	f6
	f7
	f8
	f9
	f10
	f11
	f12
	print_screen
	scroll_lock
	pause
	insert
	home
	page_up
	end
	page_down
	right
	left
	down
	up
	num_lock_clear
	kp_divide
	kp_multiply
	kp_minus
	kp_plus
	kp_enter
	kp1
	kp2
	kp3
	kp4
	kp5
	kp6
	kp7
	kp8
	kp9
	kp0
	kp_period
	application
	power
	kp_equals
	f13
	f14
	f15
	f16
	f17
	f18
	f19
	f20
	f21
	f22
	f23
	f24
	f25
	execute
	help
	menu
	@select // 'select' is a reserved keyword
	stop
	again
	undo
	cut
	copy
	paste
	find
	mute
	volume_up
	volume_down
	kp_comma
	kp_equals_as400
	alt_erase
	sys_req
	cancel
	clear
	prior
	return2
	separator
	out
	oper
	clear_again
	cr_sel
	ex_sel
	kp00
	kp000
	thousands_separator
	decimal_separator
	currency_unit
	currency_sub_unit
	kp_left_paren
	kp_right_paren
	kp_left_brace
	kp_right_brace
	kp_tab
	kp_backspace
	kp_a
	kp_b
	kp_c
	kp_d
	kp_e
	kp_f
	kp_xor
	kp_power
	kp_percent
	kp_less
	kp_greater
	kp_ampersand
	kp_dbl_ampersand
	kp_vertical_bar
	kp_dbl_vertical_bar
	kp_colon
	kp_hash
	kp_space
	kp_at
	kp_exclam
	kp_mem_store
	kp_mem_recall
	kp_mem_clear
	kp_mem_add
	kp_mem_subtract
	kp_mem_multiply
	kp_mem_divide
	kp_plus_minus
	kp_clear
	kp_clear_entry
	kp_binary
	kp_octal
	kp_decimal
	kp_hexadecimal
	l_ctrl
	l_shift
	l_alt
	l_gui
	r_ctrl
	r_shift
	r_alt
	r_gui
	mode
	sleep
	wake
	channel_increment
	channel_decrement
	media_play
	media_pause
	media_record
	media_fast_forward
	media_rewind
	media_next_track
	media_previous_track
	media_stop
	media_eject
	media_play_pause
	media_select
	ac_new
	ac_open
	ac_close
	ac_exit
	ac_save
	ac_print
	ac_properties
	ac_search
	ac_home
	ac_back
	ac_forward
	ac_stop
	ac_refresh
	ac_bookmarks
	soft_left
	soft_right
	call
	end_call
	left_tab
	level5_shift
	multi_key_compose
	l_meta
	r_meta
	l_hyper
	r_hyper
	extended_mask
	scancode_mask
}